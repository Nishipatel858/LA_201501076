`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//Name    : Nishi Patel(BTech-ICT ,sem 3)
//Subject : LA Assignment
//Topic 	 : To find inverse of a matrix
//Date 	 : 7/10/2016
//Roll no : 201501076
//////////////////////////////////////////////////////////////////////////////////

module inverse_matrix(clk);

input clk;
real A[0:4][0:9];

always@(posedge clk)
begin

		A[0][0]=16'd1;
		A[0][1]=16'd2;
		A[0][2]=16'd1;
		A[0][3]=16'd0;
		A[0][4]=16'd0;
		A[0][5]=16'd1;
		A[0][6]=16'd0;
		A[0][7]=16'd0;
		A[0][8]=16'd0;
		A[0][9]=16'd0;
		
		A[1][0]=16'd0;
	   A[1][1]=16'd1;
      A[1][2]=16'd2;
      A[1][3]=16'd1;
      A[1][4]=16'd0;
		A[1][5]=16'd0;
		A[1][6]=16'd1;
		A[1][7]=16'd0;
		A[1][8]=16'd0;
		A[1][9]=16'd0;

		A[2][0]=16'd0;
      A[2][1]=16'd0;
		A[2][2]=16'd1;
		A[2][3]=16'd2;
		A[2][4]=16'd1;
		A[2][5]=16'd0;
		A[2][6]=16'd0;
		A[2][7]=16'd1;
		A[2][8]=16'd0;
		A[2][9]=16'd0;
		
		
		A[3][0]=16'd0;
		A[3][1]=16'd0;
		A[3][2]=16'd0;
		A[3][3]=16'd1;
		A[3][4]=16'd2;
		A[3][5]=16'd0;
		A[3][6]=16'd0;
		A[3][7]=16'd0;
		A[3][8]=16'd1;
		A[3][9]=16'd0;
		
		A[4][0]=16'd0;
		A[4][1]=16'd0;
		A[4][2]=16'd0;
		A[4][3]=16'd0;
		A[4][4]=16'd1;
		A[4][5]=16'd0;
		A[4][6]=16'd0;
		A[4][7]=16'd0;
		A[4][8]=16'd0;
		A[4][9]=16'd1;


		if(A[0][0]!=0)
		begin
		A[0][0]=A[0][0]/A[0][0];
		A[0][1]=A[0][1]/A[0][0];
		A[0][2]=A[0][2]/A[0][0];
		A[0][3]=A[0][3]/A[0][0];
		A[0][4]=A[0][4]/A[0][0];
		A[0][5]=A[0][5]/A[0][0];
		A[0][6]=A[0][6]/A[0][0];
		A[0][7]=A[0][7]/A[0][0];
		A[0][8]=A[0][8]/A[0][0];
		A[0][9]=A[0][9]/A[0][0];
		
		A[1][0]=A[1][0]+(-A[1][0]*A[0][0]);
		A[1][1]=A[1][1]+(-A[1][0]*A[0][1]);
		A[1][2]=A[1][2]+(-A[1][0]*A[0][2]);
		A[1][3]=A[1][3]+(-A[1][0]*A[0][3]);
		A[1][4]=A[1][4]+(-A[1][0]*A[0][4]);
		A[1][5]=A[1][5]+(-A[1][0]*A[0][5]);
		A[1][6]=A[1][6]+(-A[1][0]*A[0][6]);
		A[1][7]=A[1][7]+(-A[1][0]*A[0][7]);
		A[1][8]=A[1][8]+(-A[1][0]*A[0][8]);
		A[1][9]=A[1][9]+(-A[1][0]*A[0][9]);
		
		
		
		
		A[2][0]=A[2][0]+(-A[2][0]*A[0][0]);
		A[2][1]=A[2][1]+(-A[2][0]*A[0][1]);
		A[2][2]=A[2][2]+(-A[2][0]*A[0][2]);
		A[2][3]=A[2][3]+(-A[2][0]*A[0][3]);
		A[2][4]=A[2][4]+(-A[2][0]*A[0][4]);
		A[2][5]=A[2][5]+(-A[2][0]*A[0][5]);
		A[2][6]=A[2][6]+(-A[2][0]*A[0][6]);
		A[2][7]=A[2][7]+(-A[2][0]*A[0][7]);
		A[2][8]=A[2][8]+(-A[2][0]*A[0][8]);
		A[2][9]=A[2][9]+(-A[2][0]*A[0][9]);
		
				
		
		A[3][0]=A[3][0]+(-A[3][0]*A[0][0]);
		A[3][1]=A[3][1]+(-A[3][0]*A[0][1]);
		A[3][2]=A[3][2]+(-A[3][0]*A[0][2]);
		A[3][3]=A[3][3]+(-A[3][0]*A[0][3]);
		A[3][4]=A[3][4]+(-A[3][0]*A[0][4]);
		A[3][5]=A[3][5]+(-A[3][0]*A[0][5]);
		A[3][6]=A[3][6]+(-A[3][0]*A[0][6]);
		A[3][7]=A[3][7]+(-A[3][0]*A[0][7]);
		A[3][8]=A[3][8]+(-A[3][0]*A[0][8]);
		A[3][9]=A[3][9]+(-A[3][0]*A[0][9]);

				
		
		A[4][0]=A[4][0]+(-A[4][0]*A[0][0]);
		A[4][1]=A[4][1]+(-A[4][0]*A[0][1]);
		A[4][2]=A[4][2]+(-A[4][0]*A[0][2]);
		A[4][3]=A[4][3]+(-A[4][0]*A[0][3]);
		A[4][4]=A[4][4]+(-A[4][0]*A[0][4]);
		A[4][5]=A[4][5]+(-A[4][0]*A[0][5]);
		A[4][6]=A[4][6]+(-A[4][0]*A[0][6]);
		A[4][7]=A[4][7]+(-A[4][0]*A[0][7]);
		A[4][8]=A[4][8]+(-A[4][0]*A[0][8]);
		A[4][9]=A[4][9]+(-A[4][0]*A[0][9]);

		end
		if(A[1][1]!=0)
		begin
		A[1][0]=A[1][0]/A[1][1];
		A[1][1]=A[1][1]/A[1][1];
		A[1][2]=A[1][2]/A[1][1];
		A[1][3]=A[1][3]/A[1][1];
		A[1][4]=A[1][4]/A[1][1];
		A[1][5]=A[1][5]/A[1][1];
		A[1][6]=A[1][6]/A[1][1];
		A[1][7]=A[1][7]/A[1][1];
		A[1][8]=A[1][8]/A[1][1];
		A[1][9]=A[1][9]/A[1][1];
		
		A[2][0]=A[2][0]+(-A[2][1]*A[1][0]);
		A[2][1]=A[2][1]+(-A[2][1]*A[1][1]);
		A[2][2]=A[2][2]+(-A[2][1]*A[1][2]);
		A[2][3]=A[2][3]+(-A[2][1]*A[1][3]);
		A[2][4]=A[2][4]+(-A[2][1]*A[1][4]);
		A[2][5]=A[2][5]+(-A[2][1]*A[1][5]);
		A[2][6]=A[2][6]+(-A[2][1]*A[1][6]);
		A[2][7]=A[2][7]+(-A[2][1]*A[1][7]);
		A[2][8]=A[2][8]+(-A[2][1]*A[1][8]);
		A[2][9]=A[2][9]+(-A[2][1]*A[1][9]);
		
		A[3][0]=A[3][0]+(-A[3][1]*A[1][0]);
		A[3][1]=A[3][1]+(-A[3][1]*A[1][1]);
		A[3][2]=A[3][2]+(-A[3][1]*A[1][2]);
		A[3][3]=A[3][3]+(-A[3][1]*A[1][3]);
		A[3][4]=A[3][4]+(-A[3][1]*A[1][4]);
		A[3][5]=A[3][5]+(-A[3][1]*A[1][5]);
		A[3][6]=A[3][6]+(-A[3][1]*A[1][6]);
		A[3][7]=A[3][7]+(-A[3][1]*A[1][7]);
		A[3][8]=A[3][8]+(-A[3][1]*A[1][8]);
		A[3][9]=A[3][9]+(-A[3][1]*A[1][9]);
	
		A[4][0]=A[4][0]+(-A[4][1]*A[1][0]);
		A[4][1]=A[4][1]+(-A[4][1]*A[1][1]);
		A[4][2]=A[4][2]+(-A[4][1]*A[1][2]);
		A[4][3]=A[4][3]+(-A[4][1]*A[1][3]);
		A[4][4]=A[4][4]+(-A[4][1]*A[1][4]);
		A[4][5]=A[4][5]+(-A[4][1]*A[1][5]);
		A[4][6]=A[4][6]+(-A[4][1]*A[1][6]);
		A[4][7]=A[4][7]+(-A[4][1]*A[1][7]);
		A[4][8]=A[4][8]+(-A[4][1]*A[1][8]);
		A[4][9]=A[4][9]+(-A[4][1]*A[1][9]);
		end
		if(A[2][2]!=0)
		begin
		A[2][0]=A[2][0]/A[2][2];
		A[2][1]=A[2][1]/A[2][2];
		A[2][2]=A[2][2]/A[2][2];
		A[2][3]=A[2][3]/A[2][2];
		A[2][4]=A[2][4]/A[2][2];
		A[2][5]=A[2][5]/A[2][2];
		A[2][6]=A[2][6]/A[2][2];
		A[2][7]=A[2][7]/A[2][2];
		A[2][8]=A[2][8]/A[2][2];
		A[2][9]=A[2][9]/A[2][2];
		
		A[3][0]=A[3][0]+(-A[3][2]*A[2][0]);
		A[3][1]=A[3][1]+(-A[3][2]*A[2][1]);
		A[3][2]=A[3][2]+(-A[3][2]*A[2][2]);
		A[3][3]=A[3][3]+(-A[3][2]*A[2][3]);
		A[3][4]=A[3][4]+(-A[3][2]*A[2][4]);
		A[3][5]=A[3][5]+(-A[3][2]*A[2][5]);
		A[3][6]=A[3][6]+(-A[3][2]*A[2][6]);
		A[3][7]=A[3][7]+(-A[3][2]*A[2][7]);
		A[3][8]=A[3][8]+(-A[3][2]*A[2][8]);
		A[3][9]=A[3][9]+(-A[3][2]*A[2][9]);
		
		A[4][0]=A[4][0]+(-A[4][2]*A[2][0]);
		A[4][1]=A[4][1]+(-A[4][2]*A[2][1]);
		A[4][2]=A[4][2]+(-A[4][2]*A[2][2]);
		A[4][3]=A[4][3]+(-A[4][2]*A[2][3]);
		A[4][4]=A[4][4]+(-A[4][2]*A[2][4]);
		A[4][5]=A[4][5]+(-A[4][2]*A[2][5]);
		A[4][6]=A[4][6]+(-A[4][2]*A[2][6]);
		A[4][7]=A[4][7]+(-A[4][2]*A[2][7]);
		A[4][8]=A[4][8]+(-A[4][2]*A[2][8]);
		A[4][9]=A[4][9]+(-A[4][2]*A[2][9]);
		end
		
		if(A[3][3]!=0)
		begin
		A[3][0]=A[3][0]/A[3][3];
		A[3][1]=A[3][1]/A[3][3];
		A[3][2]=A[3][2]/A[3][3];
		A[3][3]=A[3][3]/A[3][3];
		A[3][4]=A[3][4]/A[3][3];
		A[3][5]=A[3][5]/A[3][3];
		A[3][6]=A[3][6]/A[3][3];
		A[3][7]=A[3][7]/A[3][3];
		A[3][8]=A[3][8]/A[3][3];
		A[3][9]=A[3][9]/A[3][3];
		
		A[4][0]=A[4][0]+(-A[4][3]*A[3][0]);
		A[4][1]=A[4][1]+(-A[4][3]*A[3][1]);
		A[4][2]=A[4][2]+(-A[4][3]*A[3][2]);
		A[4][3]=A[4][3]+(-A[4][3]*A[3][3]);
		A[4][4]=A[4][4]+(-A[4][3]*A[3][4]);
		A[4][5]=A[4][5]+(-A[4][3]*A[3][5]);
		A[4][6]=A[4][6]+(-A[4][3]*A[3][6]);
		A[4][7]=A[4][7]+(-A[4][3]*A[3][7]);
		A[4][8]=A[4][8]+(-A[4][3]*A[3][8]);
		A[4][9]=A[4][9]+(-A[4][3]*A[3][9]);
		end
		if(A[4][4]!=0)
		begin
		A[4][0]=A[4][0]/A[4][4];
		A[4][1]=A[4][1]/A[4][4];
		A[4][2]=A[4][2]/A[4][4];
		A[4][3]=A[4][3]/A[4][4];
		A[4][4]=A[4][4]/A[4][4];
		A[4][5]=A[4][5]/A[4][4];
		A[4][6]=A[4][6]/A[4][4];
		A[4][7]=A[4][7]/A[4][4];
		A[4][8]=A[4][8]/A[4][4];
		A[4][9]=A[4][9]/A[4][4];
		end
		
		
		A[0][0]=A[0][0]+(-A[0][1]*A[1][0]);
		A[0][1]=A[0][1]+(-A[0][1]*A[1][1]);
		A[0][2]=A[0][2]+(-A[0][1]*A[1][2]);
		A[0][3]=A[0][3]+(-A[0][1]*A[1][3]);
		A[0][4]=A[0][4]+(-A[0][1]*A[1][4]);
		A[0][5]=A[0][5]+(-A[0][1]*A[1][5]);
		A[0][6]=A[0][6]+(-A[0][1]*A[1][6]);
		A[0][7]=A[0][7]+(-A[0][1]*A[1][7]);
		A[0][8]=A[0][8]+(-A[0][1]*A[1][8]);
		A[0][9]=A[0][9]+(-A[0][1]*A[1][9]);
		
		A[1][0]=A[1][0]+(-A[1][2]*A[2][0]);
		A[1][1]=A[1][1]+(-A[1][2]*A[2][1]);
		A[1][2]=A[1][2]+(-A[1][2]*A[2][2]);
		A[1][3]=A[1][3]+(-A[1][2]*A[2][3]);
		A[1][4]=A[1][4]+(-A[1][2]*A[2][4]);
		A[1][5]=A[1][5]+(-A[1][2]*A[2][5]);
		A[1][6]=A[1][6]+(-A[1][2]*A[2][6]);
		A[1][7]=A[1][7]+(-A[1][2]*A[2][7]);
		A[1][8]=A[1][8]+(-A[1][2]*A[2][8]);
		A[1][9]=A[1][9]+(-A[1][2]*A[2][9]);
		
		A[0][0]=A[0][0]+(-A[0][2]*A[2][0]);
		A[0][1]=A[0][1]+(-A[0][2]*A[2][1]);
		A[0][2]=A[0][2]+(-A[0][2]*A[2][2]);
		A[0][3]=A[0][3]+(-A[0][2]*A[2][3]);
		A[0][4]=A[0][4]+(-A[0][2]*A[2][4]);
		A[0][5]=A[0][5]+(-A[0][2]*A[2][5]);
		A[0][6]=A[0][6]+(-A[0][2]*A[2][6]);
		A[0][7]=A[0][7]+(-A[0][2]*A[2][7]);
		A[0][8]=A[0][8]+(-A[0][2]*A[2][8]);
		A[0][9]=A[0][9]+(-A[0][2]*A[2][9]);
		
		
		A[0][0]=A[0][0]+(-A[0][3]*A[3][0]);
		A[0][1]=A[0][1]+(-A[0][3]*A[3][1]);
		A[0][2]=A[0][2]+(-A[0][3]*A[3][2]);
		A[0][3]=A[0][3]+(-A[0][3]*A[3][3]);
		A[0][4]=A[0][4]+(-A[0][3]*A[3][4]);
		A[0][5]=A[0][5]+(-A[0][3]*A[3][5]);
		A[0][6]=A[0][6]+(-A[0][3]*A[3][6]);
		A[0][7]=A[0][7]+(-A[0][3]*A[3][7]);
		A[0][8]=A[0][8]+(-A[0][3]*A[3][8]);
		A[0][9]=A[0][9]+(-A[0][3]*A[3][9]);
		
		A[1][0]=A[1][0]+(-A[1][3]*A[3][0]);
		A[1][1]=A[1][1]+(-A[1][3]*A[3][1]);
		A[1][2]=A[1][2]+(-A[1][3]*A[3][2]);
		A[1][3]=A[1][3]+(-A[1][3]*A[3][3]);
		A[1][4]=A[1][4]+(-A[1][3]*A[3][4]);
		A[1][5]=A[1][5]+(-A[1][3]*A[3][5]);
		A[1][6]=A[1][6]+(-A[1][3]*A[3][6]);
		A[1][7]=A[1][7]+(-A[1][3]*A[3][7]);
		A[1][8]=A[1][8]+(-A[1][3]*A[3][8]);
		A[1][9]=A[1][9]+(-A[1][3]*A[3][9]);
		
		A[2][0]=A[2][0]+(-A[2][3]*A[3][0]);
		A[2][1]=A[2][1]+(-A[2][3]*A[3][1]);
		A[2][2]=A[2][2]+(-A[2][3]*A[3][2]);
		A[2][3]=A[2][3]+(-A[2][3]*A[3][3]);
		A[2][4]=A[2][4]+(-A[2][3]*A[3][4]);
		A[2][5]=A[2][5]+(-A[2][3]*A[3][5]);
		A[2][6]=A[2][6]+(-A[2][3]*A[3][6]);
		A[2][7]=A[2][7]+(-A[2][3]*A[3][7]);
		A[2][8]=A[2][8]+(-A[2][3]*A[3][8]);
		A[2][9]=A[2][9]+(-A[2][3]*A[3][9]);
		
		
		
		A[0][0]=A[0][0]+(-A[0][4]*A[4][0]);
		A[0][1]=A[0][1]+(-A[0][4]*A[4][1]);
		A[0][2]=A[0][2]+(-A[0][4]*A[4][2]);
		A[0][3]=A[0][3]+(-A[0][4]*A[4][3]);
		A[0][4]=A[0][4]+(-A[0][4]*A[4][4]);
		A[0][5]=A[0][5]+(-A[0][4]*A[4][5]);
		A[0][6]=A[0][6]+(-A[0][4]*A[4][6]);
		A[0][7]=A[0][7]+(-A[0][4]*A[4][7]);
		A[0][8]=A[0][8]+(-A[0][4]*A[4][8]);
		A[0][9]=A[0][9]+(-A[0][4]*A[4][9]);
		
		A[1][0]=A[1][0]+(-A[1][4]*A[4][0]);
		A[1][1]=A[1][1]+(-A[1][4]*A[4][1]);
		A[1][2]=A[1][2]+(-A[1][4]*A[4][2]);
		A[1][3]=A[1][3]+(-A[1][4]*A[4][3]);
		A[1][4]=A[1][4]+(-A[1][4]*A[4][4]);
		A[1][5]=A[1][5]+(-A[1][4]*A[4][5]);
		A[1][6]=A[1][6]+(-A[1][4]*A[4][6]);
		A[1][7]=A[1][7]+(-A[1][4]*A[4][7]);
		A[1][8]=A[1][8]+(-A[1][4]*A[4][8]);
		A[1][9]=A[1][9]+(-A[1][4]*A[4][9]);
		
		A[2][0]=A[2][0]+(-A[2][4]*A[4][0]);
		A[2][1]=A[2][1]+(-A[2][4]*A[4][1]);
		A[2][2]=A[2][2]+(-A[2][4]*A[4][2]);
		A[2][3]=A[2][3]+(-A[2][4]*A[4][3]);
		A[2][4]=A[2][4]+(-A[2][4]*A[4][4]);
		A[2][5]=A[2][5]+(-A[2][4]*A[4][5]);
		A[2][6]=A[2][6]+(-A[2][4]*A[4][6]);
		A[2][7]=A[2][7]+(-A[2][4]*A[4][7]);
		A[2][8]=A[2][8]+(-A[2][4]*A[4][8]);
		A[2][9]=A[2][9]+(-A[2][4]*A[4][9]);
		
		A[3][0]=A[3][0]+(-A[3][4]*A[4][0]);
		A[3][1]=A[3][1]+(-A[3][4]*A[4][1]);
		A[3][2]=A[3][2]+(-A[3][4]*A[4][2]);
		A[3][3]=A[3][3]+(-A[3][4]*A[4][3]);
		A[3][4]=A[3][4]+(-A[3][4]*A[4][4]);
		A[3][5]=A[3][5]+(-A[3][4]*A[4][5]);
		A[3][6]=A[3][6]+(-A[3][4]*A[4][6]);
		A[3][7]=A[3][7]+(-A[3][4]*A[4][7]);
		A[3][8]=A[3][8]+(-A[3][4]*A[4][8]);
		A[3][9]=A[3][9]+(-A[3][4]*A[4][9]);
		

		$write("%f	",A[0][5]);
		$write("%f	",A[0][6]);
		$write("%f	",A[0][7]);
		$write("%f	",A[0][8]);
		$display("%f	",A[0][9]);
		
		$write("%f	",A[1][5]);
		$write("%f	",A[1][6]);
		$write("%f	",A[1][7]);
		$write("%f	",A[1][8]);
		$display("%f	",A[1][9]);
		
		$write("%f	",A[2][5]);
		$write("%f	",A[2][6]);
		$write("%f	",A[2][7]);
		$write("%f	",A[2][8]);
		$display("%f	",A[2][9]);
		
		$write("%f	",A[3][5]);
		$write("%f	",A[3][6]);
		$write("%f	",A[3][7]);
		$write("%f	",A[3][8]);
		$display("%f	",A[3][9]);
		
		$write("%f	",A[4][5]);
		$write("%f	",A[4][6]);
		$write("%f	",A[4][7]);
		$write("%f	",A[4][8]);
		$display("%f	",A[4][9]);
		
	
end

endmodule
